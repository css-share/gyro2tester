//////////////////////////////////////////////////////////////
//                                                          //
//                     Charles Dickinson                           //
//                      copyright 2022                      //
//                    all rights reserved                   //
//   Title  : txfifo_wrap_syn.sv                              //
//   Author : Charles Dickinson                             //
//   Date   : MAR 2022                                      //
//                                                          //
//   Notes  :                                               //
//                                                          //
//   Revision : 1.0  Inital example                         //
//                                                          //
//                                                          //
//                                                          //
//////////////////////////////////////////////////////////////


`include "gyro_parameters.vh"




module txfifo_wrap_syn ;
logic clk;
/////////////////////////////////////////////////////////////////////////////
// AXI LIGHT DECLARATION FOR cpu_txfifo_axil_if 
/////////////////////////////////////////////////////////////////////////////

 axil_rw_if  #(.AW(CPU_TXFIFO_AW),
              .PROTW(CPU_TXFIFO_PROTW),
              .DW(CPU_TXFIFO_DW),
              .STRB(CPU_TXFIFO_STRB),
              .RESPLEN(CPU_TXFIFO_RESPLEN)) 
 cpu_txfifo_axil_if       ();  


/////////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////
// AXI DECLARATION FOR txfifo_axis_if 
/////////////////////////////////////////////////////////////////////////////

 axi_strm_if #(.DW(TXFIFO_STRM_DW),
               .SW(TXFIFO_STRM_SW),
               .UW(TXFIFO_STRM_UW))
               txfifo_axis_if ();  
   


/////////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////
// AXI DECLARATION FOR txfifo_bidir0_axis_if 
/////////////////////////////////////////////////////////////////////////////

 axi_strm_if #(.DW(TXFIFO_0_STRM_DW),
               .SW(TXFIFO_0_STRM_SW),
               .UW(TXFIFO_0_STRM_UW))
               txfifo_bidir0_axis_if ();  
   


/////////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////
// AXI DECLARATION FOR txfifo_bidir1_axis_if 
/////////////////////////////////////////////////////////////////////////////

 axi_strm_if #(.DW(TXFIFO_1_STRM_DW),
               .SW(TXFIFO_1_STRM_SW),
               .UW(TXFIFO_1_STRM_UW))
               txfifo_bidir1_axis_if ();  
   


/////////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////
// AXI DECLARATION FOR txfifo_bidir2_axis_if 
/////////////////////////////////////////////////////////////////////////////

 axi_strm_if #(.DW(TXFIFO_2_STRM_DW),
               .SW(TXFIFO_2_STRM_SW),
               .UW(TXFIFO_2_STRM_UW))
               txfifo_bidir2_axis_if ();  
   


/////////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////
// ---------------------------------------------------------------------------------------------//
//         _____ __  __  ____ ___  ____  ___          _        _  ____      _     ____          //
//        |_   _|\ \/ / |  __|_ _||  __ / _ \        | \      / ||  _ \    / \   |  _ \         //
//          | |   \/ /  | |_  | | | |_ | | | |        \ \ /\ / / | |_) |  / _ \  | |_) |        //
//          | |   / /\  |  _| | | |  _|| |_| |         \ V  V /  |  _ <  / ___ \ |  __/         //
//          |_|  /_/\_\ |_|  |___||_|   \___/           \_/\_/   |_| \_||_/   \_||_|            //
//                                                                                              //
// ---------------------------------------------------------------------------------------------//
  txfifo_wrap u_txfifo_wrap (
                   .cpu_txfifo_axil_if(cpu_txfifo_axil_if.consumer),
                   .txfifo_axis_if(txfifo_axis_if.consumer),
                   .txfifo_bidir0_axis_if(txfifo_bidir0_axis_if.producer),
                   .txfifo_bidir1_axis_if(txfifo_bidir1_axis_if.producer),
                   .txfifo_bidir2_axis_if(txfifo_bidir2_axis_if.producer)
                   );


endmodule


//////////////////////////////////////////////////////////////
//                     END OF FILE                          //
//////////////////////////////////////////////////////////////
