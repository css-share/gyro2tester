//////////////////////////////////////////////////////////////
//                                                          //
//                     Charles Dickinson                           //
//                      copyright 2022                      //
//                    all rights reserved                   //
//   Title  : bidir_wrap_syn.sv                              //
//   Author : Charles Dickinson                             //
//   Date   : MAR 2022                                      //
//                                                          //
//   Notes  :                                               //
//                                                          //
//   Revision : 1.0  Inital example                         //
//                                                          //
//                                                          //
//                                                          //
//////////////////////////////////////////////////////////////


`include "gyro_parameters.vh"




module bidir_wrap_syn ;
logic clk;
/////////////////////////////////////////////////////////////////////////////
// AXI LIGHT DECLARATION FOR cpu_bidir_axil_if 
/////////////////////////////////////////////////////////////////////////////

 axil_rw_if  #(.AW(CPU_BIDIR_AW),
              .PROTW(CPU_BIDIR_PROTW),
              .DW(CPU_BIDIR_DW),
              .STRB(CPU_BIDIR_STRB),
              .RESPLEN(CPU_BIDIR_RESPLEN)) 
 cpu_bidir_axil_if       ();  


/////////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////
// AXI DECLARATION FOR txfifo_bidir0_axis_if 
/////////////////////////////////////////////////////////////////////////////

 axi_strm_if #(.DW(TXFIFO_0_STRM_DW),
               .SW(TXFIFO_0_STRM_SW),
               .UW(TXFIFO_0_STRM_UW))
               txfifo_bidir0_axis_if ();  
   


/////////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////
// AXI DECLARATION FOR txfifo_bidir1_axis_if 
/////////////////////////////////////////////////////////////////////////////

 axi_strm_if #(.DW(TXFIFO_1_STRM_DW),
               .SW(TXFIFO_1_STRM_SW),
               .UW(TXFIFO_1_STRM_UW))
               txfifo_bidir1_axis_if ();  
   


/////////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////
// AXI DECLARATION FOR txfifo_bidir2_axis_if 
/////////////////////////////////////////////////////////////////////////////

 axi_strm_if #(.DW(TXFIFO_2_STRM_DW),
               .SW(TXFIFO_2_STRM_SW),
               .UW(TXFIFO_2_STRM_UW))
               txfifo_bidir2_axis_if ();  
   


/////////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////
// AXI DECLARATION FOR bidir_rxfifo_axis_if 
/////////////////////////////////////////////////////////////////////////////

 axi_strm_if #(.DW(RXFIFO_0_STRM_DW),
               .SW(RXFIFO_0_STRM_SW),
               .UW(RXFIFO_0_STRM_UW))
               bidir_rxfifo_axis_if ();  
   


/////////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////
// ---------------------------------------------------------------------------------------//
//         ____  ___  ____   ___  ____          _        _  ____      _     ____          //
//        |  _ ||_ _||  _ \ |_ _||  _ \        | \      / ||  _ \    / \   |  _ \         //
//        | |_)/ | | | | | | | | | |_) |        \ \ /\ / / | |_) |  / _ \  | |_) |        //
//        | |_)| | | | |_| | | | |  _ <          \ V  V /  |  _ <  / ___ \ |  __/         //
//        |____/|___||____/ |___||_| \_|          \_/\_/   |_| \_||_/   \_||_|            //
//                                                                                        //
// ---------------------------------------------------------------------------------------//
  bidir_wrap u_bidir_wrap (
                   .cpu_bidir_axil_if(cpu_bidir_axil_if.consumer),
                   .txfifo_bidir0_axis_if(txfifo_bidir0_axis_if.consumer),
                   .txfifo_bidir1_axis_if(txfifo_bidir1_axis_if.consumer),
                   .txfifo_bidir2_axis_if(txfifo_bidir2_axis_if.consumer),
                   .bidir_rxfifo_axis_if(bidir_rxfifo_axis_if.producer)
                   );


endmodule


//////////////////////////////////////////////////////////////
//                     END OF FILE                          //
//////////////////////////////////////////////////////////////
