// TOP LEVEL REGISTERS 

  `define NICMAC_TX_PCS_STATS                    32'h20000000
  `define NICMAC_TX_TSMAC_STATS                  32'h20000004
  `define NICMAC_TX_PCS_TDM_STATS                32'h20000008
  `define NICMAC_TX_TDM_STATS_0                  32'h2000000c
  `define NICMAC_TX_TDM_STATS_1                  32'h20000010
  `define NICMAC_TX_RESERVED                     32'h20000014
  `define TX_ADPT_NICMAC_PREAMBLE_55_32_REG      32'h20000100
  `define TX_ADPT_NICMAC_PREAMBLE_31_0_REG       32'h20000104
  `define TX_ADPT_NICMAC_PTP_CTRL_REG            32'h20000108
  `define TX_ADPT_NICMAC_FLOW_CTRL_REG           32'h2000010c
  `define TX_ADPT_CH0_CTRL_REG                   32'h20000200
  `define TX_ADPT_CH0_STATUS_REG                 32'h20000204
  `define TX_ADPT_CH0_TS_BARRIER_MSG_CTX_REG     32'h2000022c
  `define TX_ADPT_CH0_TS_BARRIER_MSG_CTX_REG_0   32'h2000022c
  `define TX_ADPT_CH0_BARRIER_CAP_DET_REG        32'h20000230
  `define TX_ADPT_CH0_BARRIER_CAP_DET_REG_0      32'h20000230
  `define TX_ADPT_CH1_CTRL_REG                   32'h20000280
  `define TX_ADPT_CH1_STATUS_REG                 32'h20000284
  `define TX_ADPT_CH1_TS_BARRIER_MSG_CTX_REG     32'h200002ac
  `define TX_ADPT_CH1_TS_BARRIER_MSG_CTX_REG_0   32'h200002ac
  `define TX_ADPT_CH1_BARRIER_CAP_DET_REG        32'h200002b0
  `define TX_ADPT_CH1_BARRIER_CAP_DET_REG_0      32'h200002b0
  `define TX_ADPT_CH2_CTRL_REG                   32'h20000300
  `define TX_ADPT_CH2_STATUS_REG                 32'h20000304
  `define TX_ADPT_CH2_TS_BARRIER_MSG_CTX_REG     32'h2000032c
  `define TX_ADPT_CH2_TS_BARRIER_MSG_CTX_REG_0   32'h2000032c
  `define TX_ADPT_CH2_BARRIER_CAP_DET_REG        32'h20000330
  `define TX_ADPT_CH2_BARRIER_CAP_DET_REG_0      32'h20000330
  `define TX_ADPT_CH3_CTRL_REG                   32'h20000380
  `define TX_ADPT_CH3_STATUS_REG                 32'h20000384
  `define TX_ADPT_CH3_TS_BARRIER_MSG_CTX_REG     32'h200003ac
  `define TX_ADPT_CH3_TS_BARRIER_MSG_CTX_REG_0   32'h200003ac
  `define TX_ADPT_CH3_BARRIER_CAP_DET_REG        32'h200003b0
  `define TX_ADPT_CH3_BARRIER_CAP_DET_REG_0      32'h200003b0
  `define TX_FABRIC_CHAN_0_CONFIG_REG            32'h20000400
  `define TX_FABRIC_CHAN_1_CONFIG_REG            32'h20000404

  `define NICMAC_RX_PCS_STATS                    32'h2001000c
  `define NICMAC_RX_PCS_BIP_ERR                  32'h20010010
  `define NICMAC_RX_TDM_BLK_LOCK                 32'h20010014
  `define NICMAC_RX_TDM_FEC_ERR                  32'h20010018
  `define NICMAC_RX_TDM_FEC_DELAY_01             32'h2001001c
  `define NICMAC_RX_TDM_FEC_DELAY_23             32'h20010020
  `define NICMAC_RX_TDM_ERR                      32'h20010024
  `define NICMAC_RX_PCS_TDM_GBX                  32'h20010028
  `define NICMAC_RX_PCS_TDM_LANE_ALIGNER         32'h2001002c
  `define NICMAC_RX_PCS_TDM_MF_ERR               32'h20010030
  `define NICMAC_RX_PCS_TDM_MF_LEN_ERR           32'h20010034
  `define NICMAC_RX_PCS_TDM_MF_REPEAT_ERR        32'h20010038
  `define NICMAC_RX_PCS_TDM_MMISALIGNED          32'h2001003c
  `define NICMAC_RX_PCS_TDM_SYNC_ERR             32'h20010040
  `define NICMAC_RX_RSFEC_TDM_STATS_DEMUXED      32'h20010044
  `define NICMAC_RX_PCS_TDM_STATS_DEMUXED        32'h20010048
  `define NICMAC_RX_TSMAC_TDM_STATS_PACKED       32'h2001004c
  `define NICMAC_RX_TSMAC_TDM_STATS_TOTALS       32'h20010050
  `define NICMAC_RX_TSMAC_TDM_STATS              32'h20010054
  `define NICMAC_RX_RESERVED                     32'h20010058
  `define NICMAC_RX_BS_PCS0                      32'h2001005c
  `define NICMAC_RX_BS_PCS1                      32'h2001005c
  `define NICMAC_RX_BS_PCS2                      32'h20010060
  `define NICMAC_RX_BS_PCS3                      32'h20010064
  `define NICMAC_RX_BS_TSMAC0                    32'h20010064
  `define NICMAC_RX_BS_TSMAC1                    32'h20010068
  `define NICMAC_RX_BS_TSMAC2                    32'h2001006c
  `define NICMAC_RX_BS_TSMAC3                    32'h20010070
  `define RX_ADPT_GLOBAL_CTRL_REG                32'h20010100
  `define RX_ADPT_ICSB_CALENDAR_CTRL_REG         32'h20010104
  `define RX_ADPT_ICSB_CALENDAR_SEQ_REG          32'h20010108
  `define RX_ADPT_CH0_CTRL_REG                   32'h20010200
  `define RX_ADPT_CH0_STATUS_REG                 32'h20010204
  `define RX_ADPT_CH1_CTRL_REG                   32'h20010280
  `define RX_ADPT_CH1_STATUS_REG                 32'h20010284
  `define RX_ADPT_CH2_CTRL_REG                   32'h20010300
  `define RX_ADPT_CH2_STATUS_REG                 32'h20010304
  `define RX_ADPT_CH3_CTRL_REG                   32'h20010380
  `define RX_ADPT_CH3_STATUS_REG                 32'h20010384
  `define RX_ADPT_FC_CTRL                        32'h20010400
  `define RX_ADPT_FC_DEST_MSG_MOD_CTRL           32'h20010404

  `define PDMA_WR_CFG_REG                        32'h20014000
  `define PDMA_RD_CFG_REG                        32'h20014004
  `define PDMA_MASK_A0_REG                       32'h20014008
  `define PDMA_MASK_A1_REG                       32'h2001400c
  `define PDMA_MASK_A2_REG                       32'h20014010
  `define PDMA_MASK_A3_REG                       32'h20014014
  `define PDMA_MASK_A4_REG                       32'h20014018
  `define PDMA_MASK_A5_REG                       32'h2001401c
  `define PDMA_MASK_B0_REG                       32'h20014020
  `define PDMA_MASK_B1_REG                       32'h20014024
  `define PDMA_MASK_B2_REG                       32'h20014028
  `define PDMA_MASK_B3_REG                       32'h2001402c
  `define PDMA_MASK_B4_REG                       32'h20014030
  `define PDMA_MASK_B5_REG                       32'h20014034
  `define PDMA_MASK_C0_REG                       32'h20014038
  `define PDMA_MASK_C1_REG                       32'h2001403c
  `define PDMA_MASK_C2_REG                       32'h20014040
  `define PDMA_MASK_C3_REG                       32'h20014044
  `define PDMA_MASK_C4_REG                       32'h20014048
  `define PDMA_MASK_C5_REG                       32'h2001404c
  `define PDMA_MASK_D0_REG                       32'h20014050
  `define PDMA_MASK_D1_REG                       32'h20014054
  `define PDMA_MASK_D2_REG                       32'h20014058
  `define PDMA_MASK_D3_REG                       32'h2001405c
  `define PDMA_MASK_D4_REG                       32'h20014060
  `define PDMA_MASK_D5_REG                       32'h20014064
  `define PDMA_MASK_E0_REG                       32'h20014068
  `define PDMA_MASK_E1_REG                       32'h2001406c
  `define PDMA_MASK_E2_REG                       32'h20014070
  `define PDMA_MASK_E3_REG                       32'h20014074
  `define PDMA_MASK_E4_REG                       32'h20014078
  `define PDMA_MASK_E5_REG                       32'h2001407c
  `define PDMA_MASK_F0_REG                       32'h20014080
  `define PDMA_MASK_F1_REG                       32'h20014084
  `define PDMA_MASK_F2_REG                       32'h20014088
  `define PDMA_MASK_F3_REG                       32'h2001408c
  `define PDMA_MASK_F4_REG                       32'h20014090
  `define PDMA_MASK_F5_REG                       32'h20014094
  `define PDMA_MASK_G0_REG                       32'h20014098
  `define PDMA_MASK_G1_REG                       32'h2001409c
  `define PDMA_MASK_G2_REG                       32'h200140a0
  `define PDMA_MASK_G3_REG                       32'h200140a4
  `define PDMA_MASK_G4_REG                       32'h200140a8
  `define PDMA_MASK_G5_REG                       32'h200140ac
  `define PDMA_MASK_H0_REG                       32'h200140b0
  `define PDMA_MASK_H1_REG                       32'h200140b4
  `define PDMA_MASK_H2_REG                       32'h200140b8
  `define PDMA_MASK_H3_REG                       32'h200140bc
  `define PDMA_MASK_H4_REG                       32'h200140c0
  `define PDMA_MASK_H5_REG                       32'h200140c4
  `define PDMA_MATCH_A0_REG                      32'h20014108
  `define PDMA_MATCH_A1_REG                      32'h2001410c
  `define PDMA_MATCH_A2_REG                      32'h20014110
  `define PDMA_MATCH_A3_REG                      32'h20014114
  `define PDMA_MATCH_A4_REG                      32'h20014118
  `define PDMA_MATCH_A5_REG                      32'h2001411c
  `define PDMA_MATCH_B0_REG                      32'h20014120
  `define PDMA_MATCH_B1_REG                      32'h20014124
  `define PDMA_MATCH_B2_REG                      32'h20014128
  `define PDMA_MATCH_B3_REG                      32'h2001412c
  `define PDMA_MATCH_B4_REG                      32'h20014130
  `define PDMA_MATCH_B5_REG                      32'h20014134
  `define PDMA_MATCH_C0_REG                      32'h20014138
  `define PDMA_MATCH_C1_REG                      32'h2001413c
  `define PDMA_MATCH_C2_REG                      32'h20014140
  `define PDMA_MATCH_C3_REG                      32'h20014144
  `define PDMA_MATCH_C4_REG                      32'h20014148
  `define PDMA_MATCH_C5_REG                      32'h2001414c
  `define PDMA_MATCH_D0_REG                      32'h20014150
  `define PDMA_MATCH_D1_REG                      32'h20014154
  `define PDMA_MATCH_D2_REG                      32'h20014158
  `define PDMA_MATCH_D3_REG                      32'h2001415c
  `define PDMA_MATCH_D4_REG                      32'h20014160
  `define PDMA_MATCH_D5_REG                      32'h20014164
  `define PDMA_MATCH_E0_REG                      32'h20014168
  `define PDMA_MATCH_E1_REG                      32'h2001416c
  `define PDMA_MATCH_E2_REG                      32'h20014170
  `define PDMA_MATCH_E3_REG                      32'h20014174
  `define PDMA_MATCH_E4_REG                      32'h20014178
  `define PDMA_MATCH_E5_REG                      32'h2001417c
  `define PDMA_MATCH_F0_REG                      32'h20014180
  `define PDMA_MATCH_F1_REG                      32'h20014184
  `define PDMA_MATCH_F2_REG                      32'h20014188
  `define PDMA_MATCH_F3_REG                      32'h2001418c
  `define PDMA_MATCH_F4_REG                      32'h20014190
  `define PDMA_MATCH_F5_REG                      32'h20014194
  `define PDMA_MATCH_G0_REG                      32'h20014198
  `define PDMA_MATCH_G1_REG                      32'h2001419c
  `define PDMA_MATCH_G2_REG                      32'h200141a0
  `define PDMA_MATCH_G3_REG                      32'h200141a4
  `define PDMA_MATCH_G4_REG                      32'h200141a8
  `define PDMA_MATCH_G5_REG                      32'h200141ac
  `define PDMA_MATCH_H0_REG                      32'h200141b0
  `define PDMA_MATCH_H1_REG                      32'h200141b4
  `define PDMA_MATCH_H2_REG                      32'h200141b8
  `define PDMA_MATCH_H3_REG                      32'h200141bc
  `define PDMA_MATCH_H4_REG                      32'h200141c0
  `define PDMA_MATCH_H5_REG                      32'h200141c4
  `define PDMA_PSEUDOHEAD_A0_REG                 32'h20014200
  `define PDMA_PSEUDOHEAD_A1_REG                 32'h20014204
  `define PDMA_PSEUDOHEAD_A2_REG                 32'h20014208
  `define PDMA_PSEUDOHEAD_A3_REG                 32'h2001420c
  `define PDMA_PSEUDOHEAD_A4_REG                 32'h20014210
  `define PDMA_PSEUDOHEAD_A5_REG                 32'h20014214
  `define PDMA_PSEUDOHEAD_A6_REG                 32'h20014218
  `define PDMA_PSEUDOHEAD_B0_REG                 32'h2001421c
  `define PDMA_PSEUDOHEAD_B1_REG                 32'h20014220
  `define PDMA_PSEUDOHEAD_B2_REG                 32'h20014224
  `define PDMA_PSEUDOHEAD_B3_REG                 32'h20014228
  `define PDMA_PSEUDOHEAD_B4_REG                 32'h2001422c
  `define PDMA_PSEUDOHEAD_B5_REG                 32'h20014230
  `define PDMA_PSEUDOHEAD_B6_REG                 32'h20014234


  `define PTP_CFG_ADJ_C0_REG                     32'h20018000
  `define PTP_CFG_C0_REG                         32'h20018004
  `define PTP_CFG_ADJ_C1_REG                     32'h20018008
  `define PTP_CFG_C1_REG                         32'h2001800c
  `define PTP_CFG_ADJ_C2_REG                     32'h20018010
  `define PTP_CFG_C2_REG                         32'h20018014
  `define PTP_CFG_ADJ_C3_REG                     32'h20018018
  `define PTP_CFG_C3_REG                         32'h2001801c
  `define PTP_RXDWNCNT_CH02_REG                  32'h20018020
  `define PTP_RXDWNCNT_CH35_REG                  32'h20018024
  `define PTP_TXDWNCNT_CH02_REG                  32'h20018024
  `define PTP_TXDWNCNT_CH35_REG                  32'h20018028
  `define PTP_MIPS_BUS_REG                       32'h20018080


  `define NICMAC_ID_REG                          32'h20020000
   
  `define NET_RX_REG_WA                          32'h2001C020

