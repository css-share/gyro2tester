//////////////////////////////////////////////////////////////
//                                                          //
//                     Charles Dickinson                           //
//                      copyright 2022                      //
//                    all rights reserved                   //
//   Title  : axi_inter_wrap_syn.sv                              //
//   Author : Charles Dickinson                             //
//   Date   : MAR 2022                                      //
//                                                          //
//   Notes  :                                               //
//                                                          //
//   Revision : 1.0  Inital example                         //
//                                                          //
//                                                          //
//                                                          //
//////////////////////////////////////////////////////////////


`include "gyro_parameters.vh"




module axi_inter_wrap_syn ;
logic clk;
/////////////////////////////////////////////////////////////////////////////
// AXI LIGHT DECLARATION FOR cpu_bidir_axil_if 
/////////////////////////////////////////////////////////////////////////////

 axil_rw_if  #(.AW(CPU_BIDIR_AW),
              .PROTW(CPU_BIDIR_PROTW),
              .DW(CPU_BIDIR_DW),
              .STRB(CPU_BIDIR_STRB),
              .RESPLEN(CPU_BIDIR_RESPLEN)) 
 cpu_bidir_axil_if       ();  


/////////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////
// AXI LIGHT DECLARATION FOR cpu_txfifo_axil_if 
/////////////////////////////////////////////////////////////////////////////

 axil_rw_if  #(.AW(CPU_TXFIFO_AW),
              .PROTW(CPU_TXFIFO_PROTW),
              .DW(CPU_TXFIFO_DW),
              .STRB(CPU_TXFIFO_STRB),
              .RESPLEN(CPU_TXFIFO_RESPLEN)) 
 cpu_txfifo_axil_if       ();  


/////////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////
// AXI LIGHT DECLARATION FOR cpu_rxfifo_axil_if 
/////////////////////////////////////////////////////////////////////////////

 axil_rw_if  #(.AW(CPU_RXFIFO_AW),
              .PROTW(CPU_RXFIFO_PROTW),
              .DW(CPU_RXFIFO_DW),
              .STRB(CPU_RXFIFO_STRB),
              .RESPLEN(CPU_RXFIFO_RESPLEN)) 
 cpu_rxfifo_axil_if       ();  


/////////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////
// AXI LIGHT DECLARATION FOR cpu_dma_axil_if 
/////////////////////////////////////////////////////////////////////////////

 axil_rw_if  #(.AW(CPU_DMA_AW),
              .PROTW(CPU_DMA_PROTW),
              .DW(CPU_DMA_DW),
              .STRB(CPU_DMA_STRB),
              .RESPLEN(CPU_DMA_RESPLEN)) 
 cpu_dma_axil_if       ();  


/////////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////
// AXI LIGHT DECLARATION FOR cpu_spi_axil_if 
/////////////////////////////////////////////////////////////////////////////

 axil_rw_if  #(.AW(CPU_SPI_AW),
              .PROTW(CPU_SPI_PROTW),
              .DW(CPU_SPI_DW),
              .STRB(CPU_SPI_STRB),
              .RESPLEN(CPU_SPI_RESPLEN)) 
 cpu_spi_axil_if       ();  


/////////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////
// AXI LIGHT DECLARATION FOR cpu_master_axil_if 
/////////////////////////////////////////////////////////////////////////////

 axil_rw_if  #(.AW(CPU_MASTER_AW),
              .PROTW(CPU_MASTER_PROTW),
              .DW(CPU_MASTER_DW),
              .STRB(CPU_MASTER_STRB),
              .RESPLEN(CPU_MASTER_RESPLEN)) 
 cpu_master_axil_if       ();  


/////////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////
// ---------------------------------------------------------------------------------------------------------------------//
//            _    __  __  ___         ___  _   _  _____  _____ ____          _        _  ____      _     ____          //
//           / \   \ \/ / |_ _|       |_ _|| \ | ||_   _|| ____|  _ \        | \      / ||  _ \    / \   |  _ \         //
//          / _ \   \/ /   | |         | | |  \| |  | |  |  _| | |_) |        \ \ /\ / / | |_) |  / _ \  | |_) |        //
//         / ___ \  / /\   | |         | | | |\  |  | |  | |___|  _ <          \ V  V /  |  _ <  / ___ \ |  __/         //
//        |_/   \_|/_/\_\ |___|       |___||_| \_|  |_|  |_____|_| \_|          \_/\_/   |_| \_||_/   \_||_|            //
//                                                                                                                      //
// ---------------------------------------------------------------------------------------------------------------------//
  axi_inter_wrap u_axi_inter_wrap (
                   .cpu_bidir_axil_if(cpu_bidir_axil_if.producer),
                   .cpu_txfifo_axil_if(cpu_txfifo_axil_if.producer),
                   .cpu_rxfifo_axil_if(cpu_rxfifo_axil_if.producer),
                   .cpu_dma_axil_if(cpu_dma_axil_if.producer),
                   .cpu_spi_axil_if(cpu_spi_axil_if.producer),
                   .cpu_master_axil_if(cpu_master_axil_if.consumer)
                   );


endmodule


//////////////////////////////////////////////////////////////
//                     END OF FILE                          //
//////////////////////////////////////////////////////////////
