//////////////////////////////////////////////////////////////
//                                                          //
//                     Charles Dickinson                           //
//                      copyright 2022                      //
//                    all rights reserved                   //
//   Title  : spi_1_0_wrap_syn.sv                              //
//   Author : Charles Dickinson                             //
//   Date   : MAR 2022                                      //
//                                                          //
//   Notes  :                                               //
//                                                          //
//   Revision : 1.0  Inital example                         //
//                                                          //
//                                                          //
//                                                          //
//////////////////////////////////////////////////////////////


`include "gyro_parameters.vh"




module spi_1_0_wrap_syn ;
logic clk;
/////////////////////////////////////////////////////////////////////////////
// AXI LIGHT DECLARATION FOR cpu_spi_axil_if 
/////////////////////////////////////////////////////////////////////////////

 axil_rw_if  #(.AW(CPU_SPI_AW),
              .PROTW(CPU_SPI_PROTW),
              .DW(CPU_SPI_DW),
              .STRB(CPU_SPI_STRB),
              .RESPLEN(CPU_SPI_RESPLEN)) 
 cpu_spi_axil_if       ();  


/////////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////
// ------------------------------------------------------------------------------------------------------//
//         ____   ____   ___         __           ___          _        _  ____      _     ____          //
//        / ___| |  _ \ |_ _|       /  |         / _ \        | \      / ||  _ \    / \   |  _ \         //
//        \___ \ | |_) | | |         | |        | | | |        \ \ /\ / / | |_) |  / _ \  | |_) |        //
//         ___)  |  __/  | |         | |        | |_| |         \ V  V /  |  _ <  / ___ \ |  __/         //
//        |____/ |_|    |___|        |_|         \___/           \_/\_/   |_| \_||_/   \_||_|            //
//                                                                                                       //
// ------------------------------------------------------------------------------------------------------//
  spi_1_0_wrap u_spi_1_0_wrap (
                   .cpu_spi_axil_if(cpu_spi_axil_if.consumer)
                   );


endmodule


//////////////////////////////////////////////////////////////
//                     END OF FILE                          //
//////////////////////////////////////////////////////////////
